library IEEE;
use IEEE.std_logic_1164.ALL;

entity char_location_tb is
end char_location_tb;

