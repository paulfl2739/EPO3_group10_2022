configuration vga_platforms_behaviour_cfg of vga_platforms is
   for behaviour
   end for;
end vga_platforms_behaviour_cfg;
