library IEEE;
use IEEE.std_logic_1164.ALL;

entity platform_tb is
end platform_tb;

