library IEEE;
use IEEE.std_logic_1164.ALL;

entity vhsync_tb is
end vhsync_tb;

