configuration spi_rom_behaviour_cfg of spi_rom is
   for behaviour
   end for;
end spi_rom_behaviour_cfg;
