library IEEE;
use IEEE.std_logic_1164.ALL;

entity platform_count_tb is
end platform_count_tb;

