library IEEE;
use IEEE.std_logic_1164.ALL;

entity test is
   port(clk : in  std_logic;
	random : out std_logic_vector(3 downto 0)
);
end test;

