library IEEE;
use IEEE.std_logic_1164.ALL;

entity full_register_tb is
end full_register_tb;

