configuration vhsync_behaviour_cfg of vhsync is
   for behaviour
   end for;
end vhsync_behaviour_cfg;
