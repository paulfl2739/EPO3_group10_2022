configuration integrate_structural_cfg of integrate is
   for structural
