configuration control_tb_behaviour_cfg of control_tb is
   for behaviour
      for all: control use configuration work.control_structural_cfg;
      end for;
   end for;
end control_tb_behaviour_cfg;
