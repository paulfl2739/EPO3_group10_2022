library IEEE;
use IEEE.std_logic_1164.ALL;

entity test_plat_tb is
end test_plat_tb;

