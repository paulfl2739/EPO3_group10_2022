library IEEE;
use IEEE.std_logic_1164.ALL;

entity control_tb is
end control_tb;

