configuration offset_count_behavioral_cfg of offset_count is
   for behavioral
   end for;
end offset_count_behavioral_cfg;
