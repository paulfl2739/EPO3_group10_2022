configuration char_location_behaviour_cfg of char_location is
   for behaviour
   end for;
end char_location_behaviour_cfg;
