configuration spc_clockgen_synthesised_cfg of spc_clockgen is
   for synthesised
      -- skipping dfqd1bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping aoi22d0bwp7t because it is not a local entity
      -- skipping oai32d1bwp7t because it is not a local entity
      -- skipping ckxor2d1bwp7t because it is not a local entity
      -- skipping or2d4bwp7t because it is not a local entity
      -- skipping edfkcnd0bwp7t because it is not a local entity
      -- skipping aoi21d0bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
   end for;
end spc_clockgen_synthesised_cfg;
