configuration reset_module_behavioural_cfg of reset_module is
   for behavioural
   end for;
end reset_module_behavioural_cfg;
