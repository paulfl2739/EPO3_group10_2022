configuration counter_behavioral_cfg of counter is
   for behavioral
   end for;
end counter_behavioral_cfg;
