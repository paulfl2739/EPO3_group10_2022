configuration high_edgedetec_high_edgedetector_rtl_cfg of high_edgedetec is
   for high_edgedetector_rtl
   end for;
end high_edgedetec_high_edgedetector_rtl_cfg;
