configuration clk60hz_gen_behaviour_cfg of clk60hz_gen is
   for behaviour
   end for;
end clk60hz_gen_behaviour_cfg;
