configuration top_vga_entity_structural_cfg of top_vga_entity is
   for structural
