configuration spc_clockgen_behaviour_cfg of spc_clockgen is
   for behaviour
   end for;
end spc_clockgen_behaviour_cfg;
