library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity determine_position_tb is
end entity determine_position_tb;

architecture behavioral of determine_position_tb is
    component determine_position is
        port(   clk         : in std_logic; --25 MHz internal 
        reset       : in std_logic;

        frame_passed: in std_logic; -- '1' when frame has passed for 1 clock cycle
        collision   : in std_logic; -- from VGA, duration not very important
        x_velocity   : in std_logic_vector(7 downto 0); -- from SPI

        x_position  : out std_logic_vector(8 downto 0);
        y_position  : out std_logic_vector(9 downto 0));
    end component determine_position;

    signal sig_clk, sig_reset, sig_fp, sig_col : std_logic;
    signal signedxvel : integer;
    signal sig_xvel : std_logic_vector(7 downto 0);
    signal sig_xpos : std_logic_vector(8 downto 0);
    signal sig_ypos : std_logic_vector(9 downto 0);

    begin

sig_clk <= '0' after 0 ns,
            '1' after 20 ns when sig_clk /= '1' else '0';
sig_reset <= '1' after 0 ns,
            '0' after 50 ns;
sig_fp <= '0' after 0 ns, -- 1/60 Hz officially, '1' for 1 clk cycle
                '1' after 60 ns, -- I reduced duration for simulation ease
                '0' after 80 ns,
                '1' after 120 ns,
                '0' after 140 ns,
		'1' after 200 ns,
		'0' after 220 ns,
		'1' after 300 ns,
		'0' after 320 ns;
sig_col <= '0' after 0 ns,
		'1' after 369 ns,
		'0' after 390 ns,
		'1' after 750 ns,
		'0' after 770 ns;

signedxvel <= 0 after 0 ns,
	53 after 10 ns,
	79 after 30 ns,
	20 after 50 ns,
	35 after 70 ns,
	-10 after 90 ns,
	-70 after 110 ns,
	120 after 130 ns,
	130 after 150 ns,
	-400 after 170 ns,
	0 after 190 ns;

sig_xvel <= std_logic_vector(to_signed(signedxvel, 8));

lbldp: determine_position port map(
    clk => sig_clk,
    reset => sig_reset,
    frame_passed => sig_fp,
    collision => sig_col,
    x_velocity => sig_xvel,
    x_position => sig_xpos,
    y_position => sig_ypos);


end architecture behavioral;