configuration driver_behaviour_cfg of driver is
   for behaviour
   end for;
end driver_behaviour_cfg;
