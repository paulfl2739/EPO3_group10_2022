configuration platform_behaviour_cfg of platform is
   for behaviour
   end for;
end platform_behaviour_cfg;
