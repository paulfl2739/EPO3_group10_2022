library IEEE;
use IEEE.std_logic_1164.ALL;

entity testing_tb is
end testing_tb;

