configuration edgedetector_edgedetector_rtl_cfg of edgedetector is
   for edgedetector_rtl
   end for;
end edgedetector_edgedetector_rtl_cfg;
