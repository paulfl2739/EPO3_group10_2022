configuration spi_data_ctrl_behaviour_cfg of spi_data_ctrl is
   for behaviour
   end for;
end spi_data_ctrl_behaviour_cfg;
