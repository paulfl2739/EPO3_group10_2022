library IEEE;
use IEEE.std_logic_1164.ALL;

entity galois_tb is
end galois_tb;

