use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity L3GD20H_driver is

end entity L3GD20H_driver;
